library ieee;
use ieee.std_logic_1164.all;
--generated automatically by gen_ver.py script--
package hwver_pkg is
constant c_build_date : std_logic_vector(31 downto 0) := x"12060e00";
constant c_switch_hdl_ver : std_logic_vector(31 downto 0) := x"0508ae9f";
constant c_gencores_ver : std_logic_vector(31 downto 0) := x"05118070";
constant c_wrcores_ver : std_logic_vector(31 downto 0) := x"07efeb16";
end package;
