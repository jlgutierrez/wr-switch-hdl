library ieee;
use ieee.std_logic_1164.all;

package wrsw_txtsu_pkg is

-- t_txtsu_timestamp was here, but now it's moved to wr_endpoint_pkg.
  
end wrsw_txtsu_pkg;
