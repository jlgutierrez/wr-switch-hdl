`define ADDR_RTU_GCR                   11'h0
`define RTU_GCR_G_ENA_OFFSET 0
`define RTU_GCR_G_ENA 32'h00000001
`define RTU_GCR_MFIFOTRIG_OFFSET 1
`define RTU_GCR_MFIFOTRIG 32'h00000002
`define RTU_GCR_POLY_VAL_OFFSET 8
`define RTU_GCR_POLY_VAL 32'h00ffff00
`define RTU_GCR_RTU_VERSION_OFFSET 24
`define RTU_GCR_RTU_VERSION 32'h0f000000
`define ADDR_RTU_PSR                   11'h4
`define RTU_PSR_PORT_SEL_OFFSET 0
`define RTU_PSR_PORT_SEL 32'h000000ff
`define RTU_PSR_N_PORTS_OFFSET 8
`define RTU_PSR_N_PORTS 32'h0000ff00
`define ADDR_RTU_PCR                   11'h8
`define RTU_PCR_LEARN_EN_OFFSET 0
`define RTU_PCR_LEARN_EN 32'h00000001
`define RTU_PCR_PASS_ALL_OFFSET 1
`define RTU_PCR_PASS_ALL 32'h00000002
`define RTU_PCR_PASS_BPDU_OFFSET 2
`define RTU_PCR_PASS_BPDU 32'h00000004
`define RTU_PCR_FIX_PRIO_OFFSET 3
`define RTU_PCR_FIX_PRIO 32'h00000008
`define RTU_PCR_PRIO_VAL_OFFSET 4
`define RTU_PCR_PRIO_VAL 32'h00000070
`define RTU_PCR_B_UNREC_OFFSET 7
`define RTU_PCR_B_UNREC 32'h00000080
`define ADDR_RTU_VTR1                  11'hc
`define RTU_VTR1_VID_OFFSET 0
`define RTU_VTR1_VID 32'h00000fff
`define RTU_VTR1_FID_OFFSET 12
`define RTU_VTR1_FID 32'h000ff000
`define RTU_VTR1_DROP_OFFSET 20
`define RTU_VTR1_DROP 32'h00100000
`define RTU_VTR1_HAS_PRIO_OFFSET 21
`define RTU_VTR1_HAS_PRIO 32'h00200000
`define RTU_VTR1_PRIO_OVERRIDE_OFFSET 22
`define RTU_VTR1_PRIO_OVERRIDE 32'h00400000
`define RTU_VTR1_PRIO_OFFSET 23
`define RTU_VTR1_PRIO 32'h03800000
`define RTU_VTR1_UPDATE_OFFSET 26
`define RTU_VTR1_UPDATE 32'h04000000
`define ADDR_RTU_VTR2                  11'h10
`define RTU_VTR2_PORT_MASK_OFFSET 0
`define RTU_VTR2_PORT_MASK 32'hffffffff
`define ADDR_RTU_RX_CTR                11'h14
`define RTU_RX_CTR_FF_MAC_BR_OFFSET 0
`define RTU_RX_CTR_FF_MAC_BR 32'h00000001
`define RTU_RX_CTR_FF_MAC_RANGE_OFFSET 1
`define RTU_RX_CTR_FF_MAC_RANGE 32'h00000002
`define RTU_RX_CTR_FF_MAC_SINGLE_OFFSET 2
`define RTU_RX_CTR_FF_MAC_SINGLE 32'h00000004
`define RTU_RX_CTR_FF_MAC_LL_OFFSET 3
`define RTU_RX_CTR_FF_MAC_LL 32'h00000008
`define RTU_RX_CTR_FF_MAC_PTP_OFFSET 4
`define RTU_RX_CTR_FF_MAC_PTP 32'h00000010
`define RTU_RX_CTR_MR_ENA_OFFSET 5
`define RTU_RX_CTR_MR_ENA 32'h00000020
`define RTU_RX_CTR_AT_FMATCH_TOO_SLOW_OFFSET 6
`define RTU_RX_CTR_AT_FMATCH_TOO_SLOW 32'h00000040
`define RTU_RX_CTR_PRIO_MASK_OFFSET 8
`define RTU_RX_CTR_PRIO_MASK 32'h0000ff00
`define ADDR_RTU_RX_FF_MAC_R0          11'h18
`define RTU_RX_FF_MAC_R0_LO_OFFSET 0
`define RTU_RX_FF_MAC_R0_LO 32'hffffffff
`define ADDR_RTU_RX_FF_MAC_R1          11'h1c
`define RTU_RX_FF_MAC_R1_HI_ID_OFFSET 0
`define RTU_RX_FF_MAC_R1_HI_ID 32'h0000ffff
`define RTU_RX_FF_MAC_R1_ID_OFFSET 16
`define RTU_RX_FF_MAC_R1_ID 32'h00ff0000
`define RTU_RX_FF_MAC_R1_TYPE_OFFSET 24
`define RTU_RX_FF_MAC_R1_TYPE 32'h01000000
`define RTU_RX_FF_MAC_R1_VALID_OFFSET 25
`define RTU_RX_FF_MAC_R1_VALID 32'h02000000
`define ADDR_RTU_RX_LLF                11'h20
`define RTU_RX_LLF_FF_MASK_OFFSET 0
`define RTU_RX_LLF_FF_MASK 32'hffffffff
`define ADDR_RTU_RX_MP_R0              11'h24
`define RTU_RX_MP_R0_DST_SRC_OFFSET 0
`define RTU_RX_MP_R0_DST_SRC 32'h00000001
`define RTU_RX_MP_R0_RX_TX_OFFSET 1
`define RTU_RX_MP_R0_RX_TX 32'h00000002
`define RTU_RX_MP_R0_MASK_ID_OFFSET 16
`define RTU_RX_MP_R0_MASK_ID 32'hffff0000
`define ADDR_RTU_RX_MP_R1              11'h28
`define RTU_RX_MP_R1_MASK_OFFSET 0
`define RTU_RX_MP_R1_MASK 32'hffffffff
`define ADDR_RTU_EIC_IDR               11'h40
`define RTU_EIC_IDR_NEMPTY_OFFSET 0
`define RTU_EIC_IDR_NEMPTY 32'h00000001
`define ADDR_RTU_EIC_IER               11'h44
`define RTU_EIC_IER_NEMPTY_OFFSET 0
`define RTU_EIC_IER_NEMPTY 32'h00000001
`define ADDR_RTU_EIC_IMR               11'h48
`define RTU_EIC_IMR_NEMPTY_OFFSET 0
`define RTU_EIC_IMR_NEMPTY 32'h00000001
`define ADDR_RTU_EIC_ISR               11'h4c
`define RTU_EIC_ISR_NEMPTY_OFFSET 0
`define RTU_EIC_ISR_NEMPTY 32'h00000001
`define ADDR_RTU_UFIFO_R0              11'h50
`define RTU_UFIFO_R0_DMAC_LO_OFFSET 0
`define RTU_UFIFO_R0_DMAC_LO 32'hffffffff
`define ADDR_RTU_UFIFO_R1              11'h54
`define RTU_UFIFO_R1_DMAC_HI_OFFSET 0
`define RTU_UFIFO_R1_DMAC_HI 32'h0000ffff
`define ADDR_RTU_UFIFO_R2              11'h58
`define RTU_UFIFO_R2_SMAC_LO_OFFSET 0
`define RTU_UFIFO_R2_SMAC_LO 32'hffffffff
`define ADDR_RTU_UFIFO_R3              11'h5c
`define RTU_UFIFO_R3_SMAC_HI_OFFSET 0
`define RTU_UFIFO_R3_SMAC_HI 32'h0000ffff
`define ADDR_RTU_UFIFO_R4              11'h60
`define RTU_UFIFO_R4_VID_OFFSET 0
`define RTU_UFIFO_R4_VID 32'h00000fff
`define RTU_UFIFO_R4_PRIO_OFFSET 12
`define RTU_UFIFO_R4_PRIO 32'h00007000
`define RTU_UFIFO_R4_PID_OFFSET 16
`define RTU_UFIFO_R4_PID 32'h00ff0000
`define RTU_UFIFO_R4_HAS_VID_OFFSET 24
`define RTU_UFIFO_R4_HAS_VID 32'h01000000
`define RTU_UFIFO_R4_HAS_PRIO_OFFSET 25
`define RTU_UFIFO_R4_HAS_PRIO 32'h02000000
`define ADDR_RTU_UFIFO_CSR             11'h64
`define RTU_UFIFO_CSR_EMPTY_OFFSET 17
`define RTU_UFIFO_CSR_EMPTY 32'h00020000
`define RTU_UFIFO_CSR_USEDW_OFFSET 0
`define RTU_UFIFO_CSR_USEDW 32'h0000007f
`define ADDR_RTU_MFIFO_R0              11'h68
`define RTU_MFIFO_R0_AD_SEL_OFFSET 0
`define RTU_MFIFO_R0_AD_SEL 32'h00000001
`define ADDR_RTU_MFIFO_R1              11'h6c
`define RTU_MFIFO_R1_AD_VAL_OFFSET 0
`define RTU_MFIFO_R1_AD_VAL 32'hffffffff
`define ADDR_RTU_MFIFO_CSR             11'h70
`define RTU_MFIFO_CSR_FULL_OFFSET 16
`define RTU_MFIFO_CSR_FULL 32'h00010000
`define RTU_MFIFO_CSR_EMPTY_OFFSET 17
`define RTU_MFIFO_CSR_EMPTY 32'h00020000
`define RTU_MFIFO_CSR_USEDW_OFFSET 0
`define RTU_MFIFO_CSR_USEDW 32'h0000003f
`define BASE_RTU_ARAM                  11'h400
`define SIZE_RTU_ARAM                  32'h100
