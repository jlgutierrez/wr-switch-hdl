`define ADDR_SPLL_CSR                  6'h0
`define SPLL_CSR_PER_SEL_OFFSET 0
`define SPLL_CSR_PER_SEL 32'h0000003f
`define SPLL_CSR_N_REF_OFFSET 8
`define SPLL_CSR_N_REF 32'h00003f00
`define SPLL_CSR_N_OUT_OFFSET 16
`define SPLL_CSR_N_OUT 32'h00070000
`define ADDR_SPLL_OCCR                 6'h4
`define SPLL_OCCR_OUT_EN_OFFSET 0
`define SPLL_OCCR_OUT_EN 32'h000000ff
`define SPLL_OCCR_OUT_LOCK_OFFSET 8
`define SPLL_OCCR_OUT_LOCK 32'h0000ff00
`define ADDR_SPLL_RCER                 6'h8
`define ADDR_SPLL_OCER                 6'hc
`define ADDR_SPLL_PER_HPLL             6'h10
`define SPLL_PER_HPLL_ERROR_OFFSET 0
`define SPLL_PER_HPLL_ERROR 32'h0000ffff
`define SPLL_PER_HPLL_VALID_OFFSET 16
`define SPLL_PER_HPLL_VALID 32'h00010000
`define ADDR_SPLL_DAC_HPLL             6'h14
`define ADDR_SPLL_DAC_MAIN             6'h18
`define SPLL_DAC_MAIN_VALUE_OFFSET 0
`define SPLL_DAC_MAIN_VALUE 32'h0000ffff
`define SPLL_DAC_MAIN_DAC_SEL_OFFSET 16
`define SPLL_DAC_MAIN_DAC_SEL 32'h000f0000
`define ADDR_SPLL_DEGLITCH_THR         6'h1c
`define ADDR_SPLL_EIC_IDR              6'h20
`define SPLL_EIC_IDR_TAG_OFFSET 0
`define SPLL_EIC_IDR_TAG 32'h00000001
`define ADDR_SPLL_EIC_IER              6'h24
`define SPLL_EIC_IER_TAG_OFFSET 0
`define SPLL_EIC_IER_TAG 32'h00000001
`define ADDR_SPLL_EIC_IMR              6'h28
`define SPLL_EIC_IMR_TAG_OFFSET 0
`define SPLL_EIC_IMR_TAG 32'h00000001
`define ADDR_SPLL_EIC_ISR              6'h2c
`define SPLL_EIC_ISR_TAG_OFFSET 0
`define SPLL_EIC_ISR_TAG 32'h00000001
`define ADDR_SPLL_TRR_R0               6'h30
`define SPLL_TRR_R0_VALUE_OFFSET 0
`define SPLL_TRR_R0_VALUE 32'h00ffffff
`define SPLL_TRR_R0_CHAN_ID_OFFSET 24
`define SPLL_TRR_R0_CHAN_ID 32'h7f000000
`define SPLL_TRR_R0_DISC_OFFSET 31
`define SPLL_TRR_R0_DISC 32'h80000000
`define ADDR_SPLL_TRR_CSR              6'h34
`define SPLL_TRR_CSR_EMPTY_OFFSET 17
`define SPLL_TRR_CSR_EMPTY 32'h00020000
