-------------------------------------------------------------------------------
-- Title      : multiport page allocator
-- Project    : WhiteRabbit switch
-------------------------------------------------------------------------------
-- File       : swc_multiport_page_allocator.vhd
-- Author     : Tomasz Wlostowski
-- Company    : CERN BE-Co-HT
-- Created    : 2010-04-08
-- Last update: 2010-04-08
-- Platform   : FPGA-generic
-- Standard   : VHDL'87
-------------------------------------------------------------------------------
-- Description: 
-------------------------------------------------------------------------------
-- Copyright (c) 2010 Tomasz Wlostowski
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author   Description
-- 2010-04-08  1.0      twlostow Created
-- 2010-10-11  1.1      mlipinsk comments added !!!!!
-------------------------------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.swc_swcore_pkg.all;

entity swc_multiport_page_allocator is
  port (
    rst_n_i : in std_logic;
    clk_i   : in std_logic;

    alloc_i      : in  std_logic_vector(c_swc_num_ports - 1 downto 0);
    free_i       : in  std_logic_vector(c_swc_num_ports - 1 downto 0);
    alloc_done_o : out std_logic_vector(c_swc_num_ports - 1 downto 0);
    free_done_o  : out std_logic_vector(c_swc_num_ports - 1 downto 0);

    pgaddr_free_i  : in  std_logic_vector(c_swc_num_ports * c_swc_page_addr_width - 1 downto 0);
    usecnt_i       : in  std_logic_vector(c_swc_num_ports * c_swc_usecount_width - 1 downto 0);
    pgaddr_alloc_o : out std_logic_vector(c_swc_page_addr_width-1 downto 0);

    nomem_o : out std_logic
    );

end swc_multiport_page_allocator;

architecture syn of swc_multiport_page_allocator is

  signal pg_alloc      : std_logic;
  signal pg_free       : std_logic;
  signal pg_usecnt     : std_logic_vector(c_swc_usecount_width-1 downto 0);
  signal pg_addr_alloc : std_logic_vector(c_swc_page_addr_width -1 downto 0);
  signal pg_addr_free  : std_logic_vector(c_swc_page_addr_width -1 downto 0);
  signal pg_addr_valid : std_logic;
  signal pg_idle       : std_logic;
  signal pg_done       : std_logic;
  signal pg_nomem      : std_logic;

  -- vector of requests to the Round Robin arbiter
  -- both alloc and free request
  -- the address of the bit :
  -- * representing alloc request - is even [i*2]
  -- * representing free  request - is odd  [i*2 + 1]
  signal request_vec   : std_logic_vector(c_swc_num_ports*2-1 downto 0);
  
  -- address of the request which has been granted access 
  -- to page alloation core. the LSB bit indicates the kind of
  -- operation:
  -- * '0' - even address, so alloc operation
  -- * '1' - odd  address, so free  operation
  signal request_grant : std_logic_vector(4 downto 0);

  -- used to indicate to the RR arbiter to start
  -- processing next request,
  signal request_next        : std_logic;
  
  -- indicates that the granted request is valid
  signal request_grant_valid : std_logic;

  -- the number of the port to which request has been granted
  signal in_sel              : integer range 0 to c_swc_num_ports-1;
  
  -- >????
  signal in_sel_prev         : integer range 0 to c_swc_num_ports-1;
  
  -- ??
  signal af_prev             : std_logic;

  -- indicates that an alloc has been performed successfully for the 
  -- given port. Used to prevent considering the currently process
  -- port for request to RR arbiter
  signal alloc_done_feedback : std_logic_vector(c_swc_num_ports-1 downto 0);
  

  signal alloc_done          : std_logic_vector(c_swc_num_ports-1 downto 0);

  -- indicates that an free has been performed successfully for the 
  -- given port. Used to prevent considering the currently process
  -- port for request to RR arbiter
  signal free_done_feedback  : std_logic_vector(c_swc_num_ports-1 downto 0);
  signal free_done           : std_logic_vector(c_swc_num_ports-1 downto 0);
  
begin  -- syn


  -- one allocator/deallocator for all ports
  ALLOC_CORE : swc_page_allocator
    generic map (
      g_num_pages      => c_swc_packet_mem_num_pages,
      g_page_addr_bits => c_swc_page_addr_width,
      g_use_count_bits => c_swc_usecount_width)
    port map (
      clk_i          => clk_i,
      rst_n_i        => rst_n_i,
      alloc_i        => pg_alloc,
      free_i         => pg_free,
      usecnt_i       => pg_usecnt,
      pgaddr_i       => pg_addr_free,
      pgaddr_o       => pg_addr_alloc,
      pgaddr_valid_o => pg_addr_valid,
      idle_o         => pg_idle,
      done_o         => pg_done,
      nomem_o        => pg_nomem);


  -- creating request vector with 'alloc' requests at even addresses
  -- and 'free' requests on odd addresses. The condition prevents
  -- considertion of actually processed port for the request to arbiter
  gen_request_vec : for i in 0 to c_swc_num_ports - 1 generate
    request_vec(2 * i)     <= alloc_i(i) and (not (alloc_done_feedback(i) or alloc_done(i)));
    request_vec(2 * i + 1) <= free_i(i) and (not (free_done_feedback(i) or free_done(i)));
  end generate gen_request_vec;

  -- Round Robin arbiter, quite specific for the usage, since it has the "next" 
  -- input. It is used to start processing next request well in advance, to prevent
  -- unnecessary delays
  ARB : swc_rr_arbiter
    generic map (
      g_num_ports      => c_swc_num_ports * 2,
      g_num_ports_log2 => 5)
    port map (
      clk_i         => clk_i,
      rst_n_i       => rst_n_i,
      next_i        => request_next,
      request_i     => request_vec,
      grant_o       => request_grant,
      grant_valid_o => request_grant_valid);

  -- port number to which request has been granted.
  in_sel <= to_integer(unsigned(request_grant(request_grant'length-1 downto 1)));

  -- if the granted request has even address (LSB = '0'), it means that
  -- the request was of 'alloc' type
  pg_alloc <= not request_grant(0) and request_grant_valid;

  -- if the granted request has odd address (LSB = '1'), it means that
  -- the request was of 'free' type
  pg_free  <= request_grant(0) and request_grant_valid;

  -- This is special to prevent unnecessary delays.
  -- The allocator indicates that the arbiter may start
  -- processing next request as in 2 cycles, net allocator 
  -- will finish the current job and will be ready for the next one
  request_next   <= pg_done;
  
  -- the address of the allocated page
  pgaddr_alloc_o <= pg_addr_alloc;

  -- Getting the address of the page we want to free
  pg_addr_free <= pgaddr_free_i(in_sel * c_swc_page_addr_width + c_swc_page_addr_width - 1 downto in_sel * c_swc_page_addr_width);
  
  -- getting the ouser count which should be assigned to freshly allocated page
  pg_usecnt    <= usecnt_i(in_sel * c_swc_usecount_width + c_swc_usecount_width - 1 downto in_sel * c_swc_usecount_width);

  process(clk_i, rst_n_i)
  begin
    if rising_edge(clk_i) then
      if(rst_n_i = '0') then
        alloc_done_feedback <= (others => '0');
        free_done_feedback  <= (others => '0');
      else

        -- recognizing on which port the allocation/deallocation/freeing process
        -- is about to finish. It's solely for request vector composition purpose
        for i in 0 to c_swc_num_ports-1 loop
          if(pg_done = '1' and (in_sel = i)) then
            alloc_done_feedback(i) <= not request_grant(0);
            free_done_feedback(i)  <= request_grant(0);
          else
            alloc_done_feedback(i) <= '0';
            free_done_feedback(i)  <= '0';
          end if;
        end loop;  -- i

        alloc_done <= alloc_done_feedback;
        free_done  <= free_done_feedback;
      end if;
    end if;
  end process;

  alloc_done_o <= alloc_done;
  free_done_o  <= free_done;

  
end syn;
