library ieee;
use ieee.std_logic_1164.all;

entity nport_buffer is
  
  generic (
    g_num_ports : natural)

    ;

end nport_buffer;
