`define ADDR_RTU_GCR                   16'h0
`define RTU_GCR_G_ENA_OFFSET 0
`define RTU_GCR_G_ENA 32'h00000001
`define RTU_GCR_MFIFOTRIG_OFFSET 1
`define RTU_GCR_MFIFOTRIG 32'h00000002
`define RTU_GCR_POLY_VAL_OFFSET 8
`define RTU_GCR_POLY_VAL 32'h00ffff00
`define ADDR_RTU_AGR_HCAM              16'h4
`define ADDR_RTU_PCR0                  16'h8
`define RTU_PCR0_LEARN_EN_OFFSET 0
`define RTU_PCR0_LEARN_EN 32'h00000001
`define RTU_PCR0_PASS_ALL_OFFSET 1
`define RTU_PCR0_PASS_ALL 32'h00000002
`define RTU_PCR0_PASS_BPDU_OFFSET 2
`define RTU_PCR0_PASS_BPDU 32'h00000004
`define RTU_PCR0_FIX_PRIO_OFFSET 3
`define RTU_PCR0_FIX_PRIO 32'h00000008
`define RTU_PCR0_PRIO_VAL_OFFSET 4
`define RTU_PCR0_PRIO_VAL 32'h00000070
`define RTU_PCR0_B_UNREC_OFFSET 7
`define RTU_PCR0_B_UNREC 32'h00000080
`define ADDR_RTU_PCR1                  16'hc
`define RTU_PCR1_LEARN_EN_OFFSET 0
`define RTU_PCR1_LEARN_EN 32'h00000001
`define RTU_PCR1_PASS_ALL_OFFSET 1
`define RTU_PCR1_PASS_ALL 32'h00000002
`define RTU_PCR1_PASS_BPDU_OFFSET 2
`define RTU_PCR1_PASS_BPDU 32'h00000004
`define RTU_PCR1_FIX_PRIO_OFFSET 3
`define RTU_PCR1_FIX_PRIO 32'h00000008
`define RTU_PCR1_PRIO_VAL_OFFSET 4
`define RTU_PCR1_PRIO_VAL 32'h00000070
`define RTU_PCR1_B_UNREC_OFFSET 7
`define RTU_PCR1_B_UNREC 32'h00000080
`define ADDR_RTU_PCR2                  16'h10
`define RTU_PCR2_LEARN_EN_OFFSET 0
`define RTU_PCR2_LEARN_EN 32'h00000001
`define RTU_PCR2_PASS_ALL_OFFSET 1
`define RTU_PCR2_PASS_ALL 32'h00000002
`define RTU_PCR2_PASS_BPDU_OFFSET 2
`define RTU_PCR2_PASS_BPDU 32'h00000004
`define RTU_PCR2_FIX_PRIO_OFFSET 3
`define RTU_PCR2_FIX_PRIO 32'h00000008
`define RTU_PCR2_PRIO_VAL_OFFSET 4
`define RTU_PCR2_PRIO_VAL 32'h00000070
`define RTU_PCR2_B_UNREC_OFFSET 7
`define RTU_PCR2_B_UNREC 32'h00000080
`define ADDR_RTU_PCR3                  16'h14
`define RTU_PCR3_LEARN_EN_OFFSET 0
`define RTU_PCR3_LEARN_EN 32'h00000001
`define RTU_PCR3_PASS_ALL_OFFSET 1
`define RTU_PCR3_PASS_ALL 32'h00000002
`define RTU_PCR3_PASS_BPDU_OFFSET 2
`define RTU_PCR3_PASS_BPDU 32'h00000004
`define RTU_PCR3_FIX_PRIO_OFFSET 3
`define RTU_PCR3_FIX_PRIO 32'h00000008
`define RTU_PCR3_PRIO_VAL_OFFSET 4
`define RTU_PCR3_PRIO_VAL 32'h00000070
`define RTU_PCR3_B_UNREC_OFFSET 7
`define RTU_PCR3_B_UNREC 32'h00000080
`define ADDR_RTU_PCR4                  16'h18
`define RTU_PCR4_LEARN_EN_OFFSET 0
`define RTU_PCR4_LEARN_EN 32'h00000001
`define RTU_PCR4_PASS_ALL_OFFSET 1
`define RTU_PCR4_PASS_ALL 32'h00000002
`define RTU_PCR4_PASS_BPDU_OFFSET 2
`define RTU_PCR4_PASS_BPDU 32'h00000004
`define RTU_PCR4_FIX_PRIO_OFFSET 3
`define RTU_PCR4_FIX_PRIO 32'h00000008
`define RTU_PCR4_PRIO_VAL_OFFSET 4
`define RTU_PCR4_PRIO_VAL 32'h00000070
`define RTU_PCR4_B_UNREC_OFFSET 7
`define RTU_PCR4_B_UNREC 32'h00000080
`define ADDR_RTU_PCR5                  16'h1c
`define RTU_PCR5_LEARN_EN_OFFSET 0
`define RTU_PCR5_LEARN_EN 32'h00000001
`define RTU_PCR5_PASS_ALL_OFFSET 1
`define RTU_PCR5_PASS_ALL 32'h00000002
`define RTU_PCR5_PASS_BPDU_OFFSET 2
`define RTU_PCR5_PASS_BPDU 32'h00000004
`define RTU_PCR5_FIX_PRIO_OFFSET 3
`define RTU_PCR5_FIX_PRIO 32'h00000008
`define RTU_PCR5_PRIO_VAL_OFFSET 4
`define RTU_PCR5_PRIO_VAL 32'h00000070
`define RTU_PCR5_B_UNREC_OFFSET 7
`define RTU_PCR5_B_UNREC 32'h00000080
`define ADDR_RTU_PCR6                  16'h20
`define RTU_PCR6_LEARN_EN_OFFSET 0
`define RTU_PCR6_LEARN_EN 32'h00000001
`define RTU_PCR6_PASS_ALL_OFFSET 1
`define RTU_PCR6_PASS_ALL 32'h00000002
`define RTU_PCR6_PASS_BPDU_OFFSET 2
`define RTU_PCR6_PASS_BPDU 32'h00000004
`define RTU_PCR6_FIX_PRIO_OFFSET 3
`define RTU_PCR6_FIX_PRIO 32'h00000008
`define RTU_PCR6_PRIO_VAL_OFFSET 4
`define RTU_PCR6_PRIO_VAL 32'h00000070
`define RTU_PCR6_B_UNREC_OFFSET 7
`define RTU_PCR6_B_UNREC 32'h00000080
`define ADDR_RTU_PCR7                  16'h24
`define RTU_PCR7_LEARN_EN_OFFSET 0
`define RTU_PCR7_LEARN_EN 32'h00000001
`define RTU_PCR7_PASS_ALL_OFFSET 1
`define RTU_PCR7_PASS_ALL 32'h00000002
`define RTU_PCR7_PASS_BPDU_OFFSET 2
`define RTU_PCR7_PASS_BPDU 32'h00000004
`define RTU_PCR7_FIX_PRIO_OFFSET 3
`define RTU_PCR7_FIX_PRIO 32'h00000008
`define RTU_PCR7_PRIO_VAL_OFFSET 4
`define RTU_PCR7_PRIO_VAL 32'h00000070
`define RTU_PCR7_B_UNREC_OFFSET 7
`define RTU_PCR7_B_UNREC 32'h00000080
`define ADDR_RTU_PCR8                  16'h28
`define RTU_PCR8_LEARN_EN_OFFSET 0
`define RTU_PCR8_LEARN_EN 32'h00000001
`define RTU_PCR8_PASS_ALL_OFFSET 1
`define RTU_PCR8_PASS_ALL 32'h00000002
`define RTU_PCR8_PASS_BPDU_OFFSET 2
`define RTU_PCR8_PASS_BPDU 32'h00000004
`define RTU_PCR8_FIX_PRIO_OFFSET 3
`define RTU_PCR8_FIX_PRIO 32'h00000008
`define RTU_PCR8_PRIO_VAL_OFFSET 4
`define RTU_PCR8_PRIO_VAL 32'h00000070
`define RTU_PCR8_B_UNREC_OFFSET 7
`define RTU_PCR8_B_UNREC 32'h00000080
`define ADDR_RTU_PCR9                  16'h2c
`define RTU_PCR9_LEARN_EN_OFFSET 0
`define RTU_PCR9_LEARN_EN 32'h00000001
`define RTU_PCR9_PASS_ALL_OFFSET 1
`define RTU_PCR9_PASS_ALL 32'h00000002
`define RTU_PCR9_PASS_BPDU_OFFSET 2
`define RTU_PCR9_PASS_BPDU 32'h00000004
`define RTU_PCR9_FIX_PRIO_OFFSET 3
`define RTU_PCR9_FIX_PRIO 32'h00000008
`define RTU_PCR9_PRIO_VAL_OFFSET 4
`define RTU_PCR9_PRIO_VAL 32'h00000070
`define RTU_PCR9_B_UNREC_OFFSET 7
`define RTU_PCR9_B_UNREC 32'h00000080
`define ADDR_RTU_EIC_IDR               16'h40
`define RTU_EIC_IDR_NEMPTY_OFFSET 0
`define RTU_EIC_IDR_NEMPTY 32'h00000001
`define ADDR_RTU_EIC_IER               16'h44
`define RTU_EIC_IER_NEMPTY_OFFSET 0
`define RTU_EIC_IER_NEMPTY 32'h00000001
`define ADDR_RTU_EIC_IMR               16'h48
`define RTU_EIC_IMR_NEMPTY_OFFSET 0
`define RTU_EIC_IMR_NEMPTY 32'h00000001
`define ADDR_RTU_EIC_ISR               16'h4c
`define RTU_EIC_ISR_NEMPTY_OFFSET 0
`define RTU_EIC_ISR_NEMPTY 32'h00000001
`define ADDR_RTU_UFIFO_R0              16'h50
`define RTU_UFIFO_R0_DMAC_LO_OFFSET 0
`define RTU_UFIFO_R0_DMAC_LO 32'hffffffff
`define ADDR_RTU_UFIFO_R1              16'h54
`define RTU_UFIFO_R1_DMAC_HI_OFFSET 0
`define RTU_UFIFO_R1_DMAC_HI 32'h0000ffff
`define ADDR_RTU_UFIFO_R2              16'h58
`define RTU_UFIFO_R2_SMAC_LO_OFFSET 0
`define RTU_UFIFO_R2_SMAC_LO 32'hffffffff
`define ADDR_RTU_UFIFO_R3              16'h5c
`define RTU_UFIFO_R3_SMAC_HI_OFFSET 0
`define RTU_UFIFO_R3_SMAC_HI 32'h0000ffff
`define ADDR_RTU_UFIFO_R4              16'h60
`define RTU_UFIFO_R4_VID_OFFSET 0
`define RTU_UFIFO_R4_VID 32'h00000fff
`define RTU_UFIFO_R4_PRIO_OFFSET 12
`define RTU_UFIFO_R4_PRIO 32'h00007000
`define RTU_UFIFO_R4_PID_OFFSET 16
`define RTU_UFIFO_R4_PID 32'h000f0000
`define RTU_UFIFO_R4_HAS_VID_OFFSET 20
`define RTU_UFIFO_R4_HAS_VID 32'h00100000
`define RTU_UFIFO_R4_HAS_PRIO_OFFSET 21
`define RTU_UFIFO_R4_HAS_PRIO 32'h00200000
`define ADDR_RTU_UFIFO_CSR             16'h64
`define RTU_UFIFO_CSR_EMPTY_OFFSET 17
`define RTU_UFIFO_CSR_EMPTY 32'h00020000
`define RTU_UFIFO_CSR_USEDW_OFFSET 0
`define RTU_UFIFO_CSR_USEDW 32'h0000007f
`define ADDR_RTU_MFIFO_R0              16'h68
`define RTU_MFIFO_R0_AD_SEL_OFFSET 0
`define RTU_MFIFO_R0_AD_SEL 32'h00000001
`define ADDR_RTU_MFIFO_R1              16'h6c
`define RTU_MFIFO_R1_AD_VAL_OFFSET 0
`define RTU_MFIFO_R1_AD_VAL 32'hffffffff
`define ADDR_RTU_MFIFO_CSR             16'h70
`define RTU_MFIFO_CSR_FULL_OFFSET 16
`define RTU_MFIFO_CSR_FULL 32'h00010000
`define RTU_MFIFO_CSR_EMPTY_OFFSET 17
`define RTU_MFIFO_CSR_EMPTY 32'h00020000
`define RTU_MFIFO_CSR_USEDW_OFFSET 0
`define RTU_MFIFO_CSR_USEDW 32'h0000003f
`define BASE_RTU_ARAM_MAIN             16'h4000
`define SIZE_RTU_ARAM_MAIN             32'h100
`define BASE_RTU_VLAN_TAB              16'h8000
`define SIZE_RTU_VLAN_TAB              32'h1000
