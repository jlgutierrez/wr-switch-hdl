`define ADDR_WDOG_RST_CNT              4'h0
`define ADDR_WDOG_CR                   4'h4
`define WDOG_CR_PORT_OFFSET 0
`define WDOG_CR_PORT 32'h000000ff
`define WDOG_CR_RST_OFFSET 31
`define WDOG_CR_RST 32'h80000000
`define ADDR_WDOG_ACT                  4'h8
`define ADDR_WDOG_FSM                  4'hc
`define WDOG_FSM_IB_ALLOC_OFFSET 0
`define WDOG_FSM_IB_ALLOC 32'h0000000f
`define WDOG_FSM_IB_TRANS_OFFSET 4
`define WDOG_FSM_IB_TRANS 32'h000000f0
`define WDOG_FSM_IB_RCV_OFFSET 8
`define WDOG_FSM_IB_RCV 32'h00000f00
`define WDOG_FSM_IB_LL_OFFSET 12
`define WDOG_FSM_IB_LL 32'h0000f000
`define WDOG_FSM_OB_PREP_OFFSET 16
`define WDOG_FSM_OB_PREP 32'h000f0000
`define WDOG_FSM_OB_SEND_OFFSET 20
`define WDOG_FSM_OB_SEND 32'h00f00000
`define WDOG_FSM_FREE_OFFSET 24
`define WDOG_FSM_FREE 32'h0f000000
