library ieee;
use ieee.std_logic_1164.all;
--generated automatically by gen_ver.py script--
package hwver_pkg is
constant c_build_date : std_logic_vector(31 downto 0) := x"11070d00";
constant c_switch_hdl_ver : std_logic_vector(31 downto 0) := x"0aced65b";
constant c_gencores_ver : std_logic_vector(31 downto 0) := x"04beed17";
constant c_wrcores_ver : std_logic_vector(31 downto 0) := x"00aafd08";
end package;
