-------------------------------------------------------------------------------
-- Title      : A module to snoop on PTP announce messaeges
-- Project    : White Rabbit
-------------------------------------------------------------------------------
-- File       : psu_announce_snooper.vhd
-- Author     : Maciej Lip0inski
-- Company    : CERN BE-CO-HT
-- Created    : 2015-03-17
-- Last update: 2015-03-17
-- Platform   : FPGA-generic
-- Standard   : VHDL'93
-------------------------------------------------------------------------------
-- Description: this module recognizes PTP Announce messages (over 802.3 Ethernet
-- and UDP) and extracts from them required info on the fly, i.e. sequence ID and
-- clock class)
-- useful: http://wiki.hevs.ch/uit/index.php5/Standards/Ethernet_PTP/frames
-- 
-- Where            | what      |  offset  16bit words   | value
---------------------------------------------------------------------------------------------
-- Ethernet header  | EtherType | 6 from start of header       | 0x88F7 (PTP), 0x8100 (VLAN), 0x0800 (IP), 
-- VLAN tag         | EtherType | 2 from EtherType             | 0x88F7 (PTP), 0x0800 (IP)
-- IP header v4     | ProtoType | 5 from EtherType raw/tagged  | ?? bits [7:0] = 0x11 (UDP) 
-- UDP header       | DstPort   | 7 from IPv4 ProtoType        | 0x0140 (320 -> general message)
-- PTP header       | MsgType   | 1 from EtherType raw/tagged  | [3:0]=0x2 (PTPv2) and  [11:8]=0xB (announce)
-- PTP header       | MsgType   | 3 from EtherType UDP dstPort | [3:0]=0x2 (PTPv2) and  [11:8]=0xB (announce)
-- PTP header       | PortID    |10 from MsgType               | 5 words to check 
-- PTP header       | SeqID     | 1 from PortID end            | remember
-- PTP header       | SeqID     |15 from MsgType               | remember
-- PTP Announce     | ClkClass  | 9 from SeqID                 | remember
-- 
-- 
-- TODO:
-- - check which octect of the word is IPv4 ProtoType
-- - check IHL options for IP
--   http://en.wikipedia.org/wiki/IPv4#Options
-- - check whcih octect for the word of PTP msg type
-- - 
-- 
-- 
-------------------------------------------------------------------------------
--
-- Copyright (c) 2015 CERN / BE-CO-HT
--
-- This source file is free software; you can redistribute it
-- and/or modify it under the terms of the GNU Lesser General
-- Public License as published by the Free Software Foundation;
-- either version 2.1 of the License, or (at your option) any
-- later version.
--
-- This source is distributed in the hope that it will be
-- useful, but WITHOUT ANY WARRANTY; without even the implied
-- warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR
-- PURPOSE.  See the GNU Lesser General Public License for more
-- details.
--
-- You should have received a copy of the GNU Lesser General
-- Public License along with this source; if not, download it
-- from http://www.gnu.org/licenses/lgpl-2.1.html
--
-------------------------------------------------------------------------------
-- FIXME:
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author          Description
-- 2015-03-17  1.0      mlipinsk	    Created
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.psu_pkg.all;
use work.wr_fabric_pkg.all;

entity psu_announce_snooper is
  generic(
    g_port_number   : integer := 18;
    g_snoop_mode    : t_snoop_mode := TX_SEQ_ID_MODE);
  port (
    clk_sys_i : in std_logic;
    rst_n_i   : in std_logic;

    -- interface with NIC
    snk_i                 : in  t_wrf_sink_in;
    src_i                 : in  t_wrf_source_in;
    rtu_dst_port_mask_i   : in  std_logic_vector(g_port_number-1 downto 0);
    -- internal stuff

    -- access to BRAM with stored sourceClockIdentity, needed for recognision if the
    -- announce is frmo our current parent
    ptp_source_id_addr_o  : out std_logic_vector(7  downto 0); 
    ptp_source_id_data_i  :  in std_logic_vector(15 downto 0); 

    -- vector which indicates that announce msg was detected, it indicates on which port
    -- (if tx, it says to which port the frame was being sent, if rx, it says on which port
    -- the message was received)
    rxtx_detected_mask_o  : out std_logic_vector(g_port_number-1 downto 0);

    -- indicates the snooped announce seq_id (tx)
    seq_id_o              : out std_logic_vector(15 downto 0);
    seq_id_valid_o        : out std_logic;

    -- indicates the snooped clock_class (rx)
    clock_class_o         : out std_logic_vector(15 downto 0);
    clock_class_valid_o   : out std_logic;
    
    -- config:
    ignore_rx_port_id_i      :  in std_logic
    );


end psu_announce_snooper;

architecture behavioral of psu_announce_snooper is

   type t_fsm_state is (
    WAIT_SOF,
    WAIT_DATA, 
    WAIT_ETHERTYPE,
    HAS_VTAG,
    WAIT_UDP_PROTO,
    WAIT_PTP_PORT,
    WAIT_MSG_TYPE,
    WAIT_SOURCE_PORT_ID,
    CHECK_SOURCE_PORT_ID,
    SEQ_ID,
    WAIT_CLOCK_CLASS,
    WAIT_OOB
    );

   signal data               : std_logic_vector(15 downto 0);
   signal addr               : std_logic_vector( 1 downto 0);
   signal stb                : std_logic;
   signal oob_valid          : std_logic;
   signal data_valid         : std_logic;
   signal word_cnt           : unsigned(7 downto 0); -- just enough of cnt to detect interestng stuff
   signal next_offset        : unsigned(7 downto 0); -- just enough of cnt to detect interestng stuff
   signal state              : t_fsm_state;
   signal cyc_d              : std_logic;
   signal ptp_source_id_addr : unsigned(7  downto 0); 
   signal port_mask          : std_logic_vector(g_port_number-1 downto 0);
   signal detect_mask        : std_logic_vector(31 downto 0); -- for port id from OOB of 5 bits

begin   
   -- data stored in "data" is being acked by snk | data cnt is incremented
   data_valid <= '1'       when (snk_i.cyc = '1' and snk_i.stb = '1' and src_i.stall = '0' and snk_i.adr="00") else '0';
   oob_valid  <= '1'       when (snk_i.cyc = '1' and snk_i.stb = '1' and src_i.stall = '0' and snk_i.adr="01") else '0';
   data       <= snk_i.dat when (snk_i.cyc = '1' and snk_i.stb = '1' and src_i.stall = '0') else (others => '0');

   process_data: process(clk_sys_i,rst_n_i)
   begin
    if rising_edge(clk_sys_i) then
      if rst_n_i = '0' then
        word_cnt   <= (others =>'0');
        cyc_d      <= '0';
      else

        cyc_d <= snk_i.cyc;

        if(snk_i.cyc = '0') then
           word_cnt   <= (others =>'0');
        elsif(data_valid = '1') then
           word_cnt <= word_cnt + 1;
        end if;

      end if;
    end if;
   end process;


   fsm: process(clk_sys_i,rst_n_i)
   begin
   
     if rising_edge(clk_sys_i) then
       if rst_n_i = '0' then
         next_offset          <= (others=>'0');
         state                <= WAIT_SOF;
         ptp_source_id_addr   <= (others=>'0');
         seq_id_o             <= (others=>'0');
         seq_id_valid_o       <= '0';
         clock_class_o        <= (others=>'0');
         clock_class_valid_o  <= '0';
         port_mask            <= (others=>'0');
         detect_mask<= (others=>'0');
         
         
       else
         case state is

           when WAIT_SOF =>

             if(cyc_d = '0' and snk_i.cyc ='1') then
               state                <= WAIT_DATA; 
               next_offset          <= (others=>'0');
               ptp_source_id_addr   <= (others=>'0');
               seq_id_o             <= (others=>'0');
               seq_id_valid_o       <=  '0';
               clock_class_o        <= (others=>'0');
               clock_class_valid_o  <=  '0';
               port_mask            <= rtu_dst_port_mask_i;
               detect_mask          <= (others=>'0');

             end if;

           when WAIT_DATA =>

             if (word_cnt = 0 and data_valid = '1') then
               state       <= WAIT_ETHERTYPE;
               next_offset <= to_unsigned(6, next_offset'length);
             end if;

           when WAIT_ETHERTYPE =>

             if(data_valid = '1' and word_cnt = next_offset) then
               if(data    = x"88F7") then -- PTP raw ethernet frame
                 state          <= WAIT_MSG_TYPE;
                 next_offset    <= next_offset + 1; -- th word
               elsif(data = x"8100") then -- VLAN tag
                 state          <= HAS_VTAG;
                 next_offset      <= next_offset + 2; 
               elsif(data = x"0800") then -- IP frame
                 state          <= WAIT_UDP_PROTO;
                 next_offset    <= next_offset + 5; 
               else
                 state          <= WAIT_SOF; -- we are done, it's not announce
               end if;
             end if;

           when HAS_VTAG =>

             if(data_valid = '1' and word_cnt = next_offset) then

               if(data = x"88F7") then -- PTP raw ethernet frame
                 state          <= WAIT_MSG_TYPE;
                 next_offset    <= next_offset + 1;
               elsif(data = x"0800") then -- IP frame
                 state          <= WAIT_UDP_PROTO;
                 next_offset    <= next_offset + 5;
               else
                 state          <= WAIT_SOF; -- we are done, it's not announce
               end if;
             end if;

           when WAIT_UDP_PROTO =>

             if(data_valid = '1' and word_cnt = next_offset) then
               if(data(7 downto 0) = x"11") then -- 17 is the UDP protocol
                 state          <= WAIT_PTP_PORT;
                 next_offset    <= next_offset + 7;
               else
                 state <= WAIT_SOF; -- we are done, it's not announce
               end if;
             end if;

           when WAIT_PTP_PORT =>

             if(data_valid = '1' and word_cnt = next_offset) then
               if(data = x"0140") then 
                 state          <= WAIT_MSG_TYPE;
                 next_offset    <= next_offset + 3;
               else
                 state          <= WAIT_SOF; -- we are done, it's not announce
               end if;
             end if;

           when WAIT_MSG_TYPE =>

             if(data_valid = '1' and word_cnt = next_offset) then
               if(data(11 downto 8) = x"B" and data(3 downto 0) = x"2") then --Announce of PTPv2
                 state          <= WAIT_SOURCE_PORT_ID;
                 next_offset    <= next_offset + 10;
               else 
                 state          <= WAIT_SOF; -- we are done, it's not announce
               end if;
             end if;

           when WAIT_SOURCE_PORT_ID => 

             if(data_valid = '1' and word_cnt = next_offset) then
               if(g_snoop_mode = TX_SEQ_ID_MODE or ignore_rx_port_id_i = '1') then 
                 state                 <= SEQ_ID;
                 next_offset           <= next_offset + 5;
               else
                 state                 <= CHECK_SOURCE_PORT_ID;
                 ptp_source_id_addr    <= ptp_source_id_addr + 1;
                 next_offset           <= next_offset + 4;
               end if;
             end if;

           when CHECK_SOURCE_PORT_ID =>

             if(data_valid = '1') then
               if(ptp_source_id_data_i = data) then
                 if(word_cnt = next_offset) then
                   state               <= SEQ_ID;
                   next_offset         <= next_offset + 1;
                 else
                   state               <= CHECK_SOURCE_PORT_ID;
                   ptp_source_id_addr  <= ptp_source_id_addr + 1;
                 end if;
               else
                 state                 <= WAIT_SOF; -- we are done, it's not announce
               end if;
             end if;

           when SEQ_ID =>

             if(data_valid = '1' and word_cnt = next_offset) then
               seq_id_o              <= data;
               seq_id_valid_o        <= '1';
               if(g_snoop_mode = RX_CLOCK_CLASS_MODE) then
                 state               <= WAIT_CLOCK_CLASS;
                 next_offset         <= next_offset + 9;
               else
                 state               <= WAIT_SOF;
                 detect_mask(g_port_number-1 downto 0)             <= port_mask;
                 detect_mask(31              downto g_port_number) <= (others =>'0');
               end if;
             end if;

           when WAIT_CLOCK_CLASS=>

             if(data_valid = '1' and word_cnt = next_offset) then
               state                 <= WAIT_OOB;
               clock_class_o         <= data;
               clock_class_valid_o   <= '1';
             end if;

           when WAIT_OOB =>

             if(oob_valid = '1') then -- 1st OOB word
               detect_mask           <= f_onehot_decode(data(4 downto 0));
               state                 <= WAIT_SOF;
             end if;

           when others => null;

         end case;
       end if;
     end if;    
   end process;

  ptp_source_id_addr_o <=std_logic_vector(ptp_source_id_addr);
  rxtx_detected_mask_o <=detect_mask(g_port_number-1 downto 0);
end behavioral;

